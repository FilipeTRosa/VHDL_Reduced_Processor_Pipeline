library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;

entity controle is
	port(
		opcode			: in std_logic;
		brEnable		: 
		ulaOp			:
		muxUlaIn1		:
		muxBrData		:
		
	);
end entity;
architecture behavior of controle is
begin




process()
begin




end process;
end behavior;